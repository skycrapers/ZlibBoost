
    .subckt OR2X2 Y B vdd vss A
M0 a_9_54# A a_2_54# vdd PMOS_VTH w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u 
M1 vdd B a_9_54# vdd PMOS_VTH w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u 
M2 Y a_2_54# vdd vdd PMOS_VTH w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u 
M3 a_2_54# A vss vss NMOS_VTH w=0.25u l=0.05u
+ ad=0p pd=0u as=0p ps=0u 
M4 vss B a_2_54# vss NMOS_VTH w=0.25u l=0.05u
+ ad=0p pd=0u as=0p ps=0u 
M5 Y a_2_54# vss vss NMOS_VTH w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u 

.ENDS