
    .subckt NOR2X1 vdd B vss Y A
M0 a_9_54# A vdd vdd PMOS_VTH w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u 
M1 Y B a_9_54# vdd PMOS_VTH w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u 
M2 Y A vss vss NMOS_VTH w=0.25u l=0.05u
+ ad=0p pd=0u as=0p ps=0u 
M3 vss B Y vss NMOS_VTH w=0.25u l=0.05u
+ ad=0p pd=0u as=0p ps=0u 

.ENDS