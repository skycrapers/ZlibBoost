
    .subckt LATCH D Q vss vdd CLK
M0 vdd CLK a_2_6# vdd PMOS_VTH w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u 
M1 a_18_74# D vdd vdd PMOS_VTH w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u 
M2 a_23_6# a_2_6# a_18_74# vdd PMOS_VTH w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u 
M3 a_35_84# CLK a_23_6# vdd PMOS_VTH w=0.25u l=0.05u
+ ad=0p pd=0u as=0p ps=0u 
M4 vdd Q a_35_84# vdd PMOS_VTH w=0.25u l=0.05u
+ ad=0p pd=0u as=0p ps=0u 
M5 vss CLK a_2_6# vss NMOS_VTH w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u 
M6 Q a_23_6# vdd vdd PMOS_VTH w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u 
M7 a_18_6# D vss vss NMOS_VTH w=0.25u l=0.05u
+ ad=0p pd=0u as=0p ps=0u 
M8 a_23_6# CLK a_18_6# vss NMOS_VTH w=0.25u l=0.05u
+ ad=0p pd=0u as=0p ps=0u 
M9 a_35_6# a_2_6# a_23_6# vss NMOS_VTH w=0.25u l=0.05u
+ ad=0p pd=0u as=0p ps=0u 
M10 vss Q a_35_6# vss NMOS_VTH w=0.25u l=0.05u
+ ad=0p pd=0u as=0p ps=0u 
M11 Q a_23_6# vss vss NMOS_VTH w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u 

.ENDS